LIBRARY 	IEEE;
USE 		IEEE.STD_LOGIC_1164.ALL;

ENTITY UNIVERSAL_SHIFT_REGISTER IS
		PORT (
					CLOCK, CLEAR, SL_IN, SR_IN : IN BIT;
					MODE 								: IN BIT_VECTOR 	 ( 1 DOWNTO 0 );
					DATA 								: IN BIT_VECTOR 	 ( 3 DOWNTO 0 );
					Q 									: INOUT BIT_VECTOR ( 3 DOWNTO 0 )
				);
END UNIVERSAL_SHIFT_REGISTER;

ARCHITECTURE BEHAVIORAL OF UNIVERSAL_SHIFT_REGISTER IS
	BEGIN
	PROCESS (CLOCK, CLEAR)
		BEGIN 							-- ASYNCHRONOUS, ACTIVE-LOW CLEAR INPUT:
			IF CLEAR = '0' THEN
				Q <= "0000" ; 			-- RISING EDGE-TRIGGERED D FLIP-FLOPS:
				
			ELSIF CLOCK'EVENT AND CLOCK = '1' THEN
				CASE MODE IS
					WHEN "00" => NULL;				 							-- "DO NOTHING" MODE: RETAIN CURRENT FLIP-FLOP OUTPUTS
					WHEN "01" => Q <= (Q SRL 1) OR (SR_IN & "000") ; 	-- SHIFT RIGHT SERIAL INPUT
					WHEN "10" => Q <= (Q SLL 1) OR ("000" & SL_IN) ; 	-- SHIFT LEFT SERIAL INPUT
					WHEN "11" => Q <= DATA ; 									-- PARALLEL (BROADSIDE) LOAD
				END CASE;
			END IF;
	END PROCESS;
END BEHAVIORAL;
