LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
 
ENTITY RIPPLECARRYADDER IS
	PORT ( 
			A 			: IN STD_LOGIC_VECTOR 	(1 DOWNTO 0);
			B 			: IN STD_LOGIC_VECTOR 	(1 DOWNTO 0);
			CIN 		: IN STD_LOGIC;
			S 			: OUT STD_LOGIC_VECTOR 	(1 DOWNTO 0);
			COUT 		: OUT STD_LOGIC
			);
	END RIPPLECARRYADDER;
 
ARCHITECTURE BEHAVIORAL OF RIPPLECARRYADDER IS
 
	COMPONENT FULLADDER
		PORT ( 
				A 		: IN STD_LOGIC;
				B 		: IN STD_LOGIC;
				CIN 	: IN STD_LOGIC;
				S 		: OUT STD_LOGIC;
				COUT 	: OUT STD_LOGIC
				);
	END COMPONENT;
 
-- INTERMEDIATE CARRY DECLARATION
SIGNAL C1		: STD_LOGIC;
 
BEGIN
 
-- PORT MAPPING FULL ADDER 4 TIMES
FA1: FULLADDER PORT MAP( A(0), B(0), CIN, S(0), C1);
FA2: FULLADDER PORT MAP( A(1), B(1), C1, S(1), COUT);

 
END BEHAVIORAL;
