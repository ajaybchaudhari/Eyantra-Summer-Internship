LIBRARY 	IEEE;
USE 		IEEE.STD_LOGIC_1164.ALL;
USE 		IEEE.NUMERIC_STD.ALL;

ENTITY FULLADDER IS
	PORT(
			A 		: IN 	STD_LOGIC;
			B 		: IN 	STD_LOGIC;
			CIN	: IN 	STD_LOGIC;
			
			S 		: OUT STD_LOGIC;
			COUT 	: OUT STD_LOGIC
			);
	END  FULLADDER;
	
	
ARCHITECTURE BEHAVIOUR OF FULLADDER IS
	BEGIN
		
			S 		<= 	A XOR B XOR CIN;
			COUT	<=		(A AND B) OR (CIN AND (A XOR B));
			

END ARCHITECTURE BEHAVIOUR;


 